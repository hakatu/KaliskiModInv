module testbench;
parameter N = 256;
  
reg [N-1:0] A;
reg [N-1:0] P;
reg start_inv;
reg clk;
reg reset_n;

wire [N-1:0] result;
wire  done_inv;

      inv U0 (
										.clk(clk),
										.reset_n(reset_n),
										.start_inv(start_inv),
										.a(A),
										.P(P),
										.done_inv(done_inv),
										.result(result)
   );
  
initial begin
clk <= 0;
forever #1 clk <= ~clk;
end

initial begin
A = 256'd6854325554222215243052392924557410287123964824515306282021023372829163033700;
P = 256'd115792089237316195423570985008687907853269984665640564039457584007908834671663;
reset_n = 0;
start_inv = 0;
#20;
A = 256'd6854325554222215243052392924557410287123964824515306282021023372829163033700;
P = 256'd115792089237316195423570985008687907853269984665640564039457584007908834671663;
reset_n = 1;
start_inv = 1;
#20;
A = 256'd6854325554222215243052392924557410287123964824515306282021023372829163033700;
P = 256'd115792089237316195423570985008687907853269984665640564039457584007908834671663;
reset_n = 1;
start_inv = 1;
/*
#10;
A = 256'd6854325554222215243052392924557410287123964824515306282021023372829163033700;
P = 256'd115792089237316195423570985008687907853269984665640564039457584007908834671663;
reset_n = 1;
start_inv = 0;
*/
	@(done_inv) begin
	A = 256'd4;
	P = 256'd115792089237316195423570985008687907853269984665640564039457584007908834671663;
	reset_n = 1;
	start_inv = 0;
	end

end
endmodule
